`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: HA_SUB

//////////////////////////////////////////////////////////////////////////////////


module HA_SUB(
    input A,
    input B,
    output Diff,
    output Borrow
    );
    
    assign Diff = A ^ B, 
           Borrow = ~A & B;  
endmodule
