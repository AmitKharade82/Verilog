`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: XNOR

//////////////////////////////////////////////////////////////////////////////////


module XNOR(
    input A,
    input B,
    output Y
    );
    assign Y = A ~^ B;
endmodule
