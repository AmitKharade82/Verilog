`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: OR

//////////////////////////////////////////////////////////////////////////////////


module OR(
    input A,
    input B,
    output Y
    );
    assign Y = A | B; 
endmodule
