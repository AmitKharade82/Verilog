`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: NOR

//////////////////////////////////////////////////////////////////////////////////


module NOR(
    input A,
    input B,
    output Y
    );
    assign Y = ~(A | B); 
endmodule
