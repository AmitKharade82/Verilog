`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: 4_1 D-MUX

//////////////////////////////////////////////////////////////////////////////////


module  DMUX(
    input IN,
    input [1:0] S,
    output [3:0] Y
    );
    assign Y[0] =  (IN & ~S[1] & ~S[0]),
           Y[1] =  (IN & ~S[1] & S[0]),
           Y[2] =  (IN & S[1] & ~S[0]),
           Y[3] =  (IN & S[1] &S[0]);
           
endmodule
