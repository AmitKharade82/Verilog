`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: XOR

//////////////////////////////////////////////////////////////////////////////////


module XOR(
    input A,
    input B,
    output Y
    );
    assign Y = A ^ B;
endmodule
