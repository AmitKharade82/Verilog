`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: HS_SUB

//////////////////////////////////////////////////////////////////////////////////


module HS_SUB(
    input A,
    input B,
    output Diff,
    output Borrow
    );
    
    assign Diff = A ^ B, 
           Borrow = ~A & B;  
endmodule
